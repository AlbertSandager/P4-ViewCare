-- megafunction wizard: %FIR Compiler II v13.1%
-- GENERATION: XML
-- LP1000.vhd

-- Generated using ACDS version 13.1 162 at 2019.05.14.11:05:34

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LP1000 is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(23 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity LP1000;

architecture rtl of LP1000 is
	component LP1000_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(23 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component LP1000_0002;

begin

	lp1000_inst : component LP1000_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of LP1000
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2019 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
-- Retrieval info: 	<generic name="filterType" value="Single Rate" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="1" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
-- Retrieval info: 	<generic name="clockRate" value="50" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="speedGrade" value="Medium" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="inputRate" value="0.008" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="inputType" value="Signed Binary" />
-- Retrieval info: 	<generic name="inputBitWidth" value="24" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="-5.953507802473751E-5,-6.135167635343702E-5,-6.317223481274333E-5,-6.499693389104716E-5,-6.682595197290053E-5,-6.865946512061758E-5,-7.049764685557237E-5,-7.234066793929237E-5,-7.418869615445064E-5,-7.604189608586106E-5,-7.79004289015743E-5,-7.976445213418295E-5,-8.163411946243434E-5,-8.35095804932554E-5,-8.539098054429423E-5,-8.72784604270788E-5,-8.917215623089688E-5,-9.10721991075013E-5,-9.297871505674132E-5,-9.48918247132236E-5,-9.681164313410566E-5,-9.873827958812245E-5,-1.0067183734594933E-4,-1.0261241347200124E-4,-1.0456009861776952E-4,-1.065149768167974E-4,-1.0847712528139286E-4,-1.1044661420117793E-4,-1.1242350654357457E-4,-1.1440785785632266E-4,-1.1639971607212963E-4,-1.1839912131554572E-4,-1.204061057121627E-4,-1.224206932002273E-4,-1.2444289934476804E-4,-1.2647273115432201E-4,-1.2851018690035904E-4,-1.3055525593948954E-4,-1.326079185385475E-4,-1.346681457026374E-4,-1.3673589900623043E-4,-1.3881113042739677E-4,-1.4089378218525974E-4,-1.4298378658075266E-4,-1.4508106584076137E-4,-1.4718553196573517E-4,-1.492970865808406E-4,-1.5141562079073928E-4,-1.5354101503806578E-4,-1.556731389656764E-4,-1.5781185128274774E-4,-1.5995699963478998E-4,-1.6210842047764885E-4,-1.6426593895556307E-4,-1.6642936878334233E-4,-1.6859851213273206E-4,-1.707731595230259E-4,-1.729530897159882E-4,-1.751380696151447E-4,-1.773278541694991E-4,-1.7952218628172918E-4,-1.8172079672091907E-4,-1.839234040398753E-4,-1.861297144970781E-4,-1.8833942198331612E-4,-1.9055220795304766E-4,-1.9276774136053326E-4,-1.949856786007816E-4,-1.9720566345534654E-4,-1.9942732704301277E-4,-2.0165028777540683E-4,-2.0387415131756386E-4,-2.060985105534836E-4,-2.083229455567016E-4,-2.1054702356590533E-4,-2.1277029896561763E-4,-2.1499231327196932E-4,-2.172125951235829E-4,-2.1943066027758476E-4,-2.2164601161076068E-4,-2.2385813912586836E-4,-2.2606651996312025E-4,-2.2827061841684395E-4,-2.304698859573269E-4,-2.326637612578528E-4,-2.3485167022692973E-4,-2.370330260457115E-4,-2.3920722921061115E-4,-2.4137366758110148E-4,-2.4353171643269812E-4,-2.456807385151158E-4,-2.478200841155872E-4,-2.499490911273343E-4,-2.520670851231749E-4,-2.541733794342482E-4,-2.562672752338433E-4,-2.583480616263057E-4,-2.604150157410026E-4,-2.624674028313193E-4,-2.645044763786608E-4,-2.66525478201431E-4,-2.6852963856895644E-4,-2.7051617632032027E-4,-2.724842989880783E-4,-2.7443320292681064E-4,-2.7636207344647806E-4,-2.782700849505394E-4,-2.8015640107878633E-4,-2.82020174854853E-4,-2.8386054883835577E-4,-2.856766552816095E-4,-2.8746761629087875E-4,-2.8923254399210543E-4,-2.909705407010634E-4,-2.9268069909788627E-4,-2.943621024059075E-4,-2.960138245747612E-4,-2.976349304676783E-4,-2.9922447605291937E-4,-3.007815085992852E-4,-3.0230506687563296E-4,-3.037941813543404E-4,-3.0524787441864803E-4,-3.066651605738095E-4,-3.080450466619849E-4,-3.093865320808018E-4,-3.1068860900551566E-4,-3.1195026261469406E-4,-3.131704713193515E-4,-3.143482069954589E-4,-3.1548243521975267E-4,-3.1657211550876086E-4,-3.1761620156097717E-4,-3.1861364150209177E-4,-3.19563378133208E-4,-3.2046434918195707E-4,-3.2131548755643383E-4,-3.22115721601865E-4,-3.2286397535993155E-4,-3.235591688306561E-4,-3.2420021823677324E-4,-3.247860362904955E-4,-3.2531553246258917E-4,-3.2578761325367155E-4,-3.2620118246764416E-4,-3.265551414871733E-4,-3.268483895511276E-4,-3.270798240338866E-4,-3.272483407264294E-4,-3.273528341191147E-4,-3.2739219768606074E-4,-3.273653241710388E-4,-3.2727110587478563E-4,-3.2710843494364805E-4,-3.268762036594662E-4,-3.2657330473060954E-4,-3.2619863158406774E-4,-3.2575107865851426E-4,-3.2522954169824546E-4,-3.246329180479088E-4,-3.2396010694792706E-4,-3.2321000983053124E-4,-3.2238153061631006E-4,-3.2147357601118576E-4,-3.2048505580373015E-4,-3.1941488316272813E-4,-3.182619749349009E-4,-3.170252519427021E-4,-3.1570363928209473E-4,-3.142960666202276E-4,-3.1280146849291723E-4,-3.1121878460185174E-4,-3.095469601114339E-4,-3.0778494594516987E-4,-3.059316990815251E-4,-3.039861828491633E-4,-3.0194736722147637E-4,-2.9981422911033533E-4,-2.9758575265896787E-4,-2.9526092953388724E-4,-2.9283875921579165E-4,-2.9031824928935014E-4,-2.8769841573179905E-4,-2.849782832002719E-4,-2.82156885317778E-4,-2.792332649577624E-4,-2.76206474527165E-4,-2.7307557624790357E-4,-2.698396424367137E-4,-2.664977557832615E-4,-2.6304900962646776E-4,-2.594925082289659E-4,-2.558273670496255E-4,-2.520527130140718E-4,-2.481676847831353E-4,-2.4417143301916003E-4,-2.4006312065010996E-4,-2.3584192313140493E-4,-2.3150702870542182E-4,-2.2705763865860155E-4,-2.2249296757609978E-4,-2.178122435939148E-4,-2.1301470864844454E-4,-2.0809961872340194E-4,-2.030662440940416E-4,-1.9791386956863696E-4,-1.92641794727154E-4,-1.872493341570665E-4,-1.8173581768626538E-4,-1.7610059061300354E-4,-1.7034301393283207E-4,-1.6446246456247804E-4,-1.5845833556061003E-4,-1.5233003634545404E-4,-1.460769929092096E-4,-1.3969864802921707E-4,-1.3319446147584584E-4,-1.2656391021704545E-4,-1.1980648861953246E-4,-1.129217086465683E-4,-1.0590910005228389E-4,-9.876821057252495E-5,-9.149860611217436E-5,-8.409987092891577E-5,-7.657160781341133E-5,-6.891343826585312E-5,-6.112500266886022E-5,-5.320596045669486E-5,-4.51559902807569E-5,-3.697479017134127E-5,-2.866207769562532E-5,-2.0217590111854238E-5,-1.1641084519710755E-5,-2.9323380068394464E-6,5.9088522085035684E-6,1.4882668638683254E-5,2.398927339183627E-5,3.322880804094929E-5,4.260139349688798E-5,5.210712988539563E-5,6.174609642807749E-5,7.151835132738339E-5,8.142393165561031E-5,9.146285324793341E-5,1.0163511059948344E-4,1.1194067676647672E-4,1.2237950327141585E-4,1.3295152001236983E-4,1.436566351763377E-4,1.544947351567141E-4,1.6546568447485863E-4,1.7656932570577505E-4,1.8780547940791477E-4,1.9917394405709842E-4,2.1067449598457418E-4,2.223068893192031E-4,2.340708559337868E-4,2.4596610539553266E-4,2.5799232492066244E-4,2.701491793331621E-4,2.82436311027678E-4,2.9485333993655577E-4,3.0739986350102424E-4,3.2007545664651776E-4,3.328796717621447E-4,3.4581203868428665E-4,3.5887206468433925E-4,3.720592344605779E-4,3.8537301013415496E-4,3.988128312492175E-4,4.1237811477713975E-4,4.2606825512486865E-4,4.3988262414737674E-4,4.5382057116420525E-4,4.6788142298010544E-4,4.820644839097579E-4,4.96369035806571E-4,5.10794338095539E-4,5.253396278101634E-4,5.400041196334158E-4,5.547870059427447E-4,5.69687456859102E-4,5.847046202999914E-4,5.998376220365209E-4,6.150855657544465E-4,6.304475331191992E-4,6.45922583844885E-4,6.61509755767235E-4,6.772080649205063E-4,6.930165056183088E-4,7.089340505383558E-4,7.249596508111086E-4,7.41092236112319E-4,7.573307147594434E-4,7.736739738119159E-4,7.901208791752656E-4,8.066702757090665E-4,8.233209873386998E-4,8.400718171709102E-4,8.569215476131493E-4,8.738689404966794E-4,8.909127372034287E-4,9.080516587965724E-4,9.25284406154831E-4,9.426096601104665E-4,9.600260815909479E-4,9.775323117642836E-4,9.951269721879936E-4,0.0010128086649616977,0.0010305759728833177,0.0010484274596088495,0.0010663616698157123,0.0010843771293696303,0.001102472345495047,0.0011206458069490362,0.0011388959841987013,0.0011572213296020273,0.0011756202775921821,0.0011940912448652296,0.0012126326305712388,0.001231242816508769,0.0012499201673227068,0.0012686630307054232,0.001287469737601248,0.0013063386024142103,0.0013252679232190468,0.0013442559819754382,0.0013633010447454527,0.0013824013619141713,0.0014015551684134727,0.0014207606839489464,0.00144001611322991,0.0014593196462025088,0.0014786694582858606,0.001498063710611228,0.0015175005502641816,0.0015369781105297375,0.001556494511140425,0.0015760478585272663,0.0015956362460736399,0.0016152577543719858,0.0016349104514833332,0.0016545923931996142,0.0016743016233087364,0.0016940361738623725,0.001713794065446446,0.0017335733074542753,0.0017533718983623375,0.0017731878260086264,0.00179301906787356,0.001812863591363419,0.0018327193540962532,0.0018525843041902507,0.0018724563805545078,0.0018923335131821783,0.0019122136234459507,0.0019320946243958294,0.0019519744210591676,0.001971850910742915,0.001991721983338051,0.0020115855216261396,0.002031439401587993,0.0020512814927143696,0.0020711096583186915,0.0020909217558517205,0.0021107156372181584,0.002130489149095115,0.0021502401332524055,0.00216996642687464,0.0021896658628850364,0.0022093362702709273,0.002228975474410903,0.0022485812974035505,0.0022681515583977247,0.0022876840739243184,0.002307176658229464,0.0023266271236091285,0.00234603328074504,0.0023653929390418994,0.0023847039069658156,0.0024039639923839223,0.002423171002905102,0.0024423227462217895,0.0024614170304527666,0.0024804516644869132,0.002499424458327856,0.0025183332234394364,0.002537175773091972,0.0025559499227092173,0.0025746534902159855,0.00259328429638637,0.002611840165192486,0.0026303189241536954,0.0026487184046862303,0.002667036442453171,0.002685270877714688,0.002703419555678523,0.002721480326850601,0.0027394510473857424,0.002757329579438388,0.0027751137915132764,0.002792801558816015,0.0028103907636034633,0.002827879295533866,0.0028452650520166783,0.0028625459385619913,0.0028797198691295094,0.0028967847664770037,0.002913738562508161,0.0029305791986197725,0.0029473046260481885,0.0029639128062149554,0.0029804017110715746,0.0029967693234433175,0.0030130136373720065,0.003029132658457702,0.0030451244041992233,0.003060986904333421,0.0030767182011731393,0.003092316349943788,0.0031077794191184515,0.003123105490751459,0.003138292660810352,0.003153339039506163,0.0031682427516219382,0.0031830019368394302,0.0031976147500638874,0.0032120793617468574,0.0032263939582069497,0.003240556741948457,0.0032545659319777906,0.003268419764117635,0.0032821164913187538,0.0032956543839693835,0.003309031730202117,0.0033222468361982496,0.0033352980264894495,0.003348183644256752,0.0033609020516267457,0.003373451629964919,0.003385830780166072,0.0033980379229417317,0.0034100714991045097,0.0034219299698493052,0.0034336118170313202,0.003445115543440783,0.0034564396730743345,0.003467582751403001,0.003478543345636684,0.003489320044985109,0.003499911460915155,0.003510316227404508,0.0035205330011915718,0.0035305604620215728,0.0035403973128887893,0.0035500422802748535,0.0035594941143830563,0.0035687515893685936,0.0035778135035647017,0.0035866786797046145,0.0035953459651392886,0.0036038142320508415,0.0036120823776616346,0.003620149324438965,0.003628014020295289,0.003635675438783951,0.003643132579290336,0.0036503844672184198,0.0036574301541726453,0.003664268718135102,0.003670899263637934,0.0036773209219309456,0.0036835328511443557,0.003689534236446657,0.003695324290197536,0.003700902252095814,0.003706267389322367,0.0037114189966779842,0.003716356396716135,0.0037210789398705924,0.0037255860045779,0.003729876997394628,0.003733951353109393,0.0037378085348496225,0.003741448034183014,0.0037448693712136736,0.0037480720946729113,0.003751055782004644,0.003753820039445428,0.0037563645020990393,0.0037586888340056354,0.0037607927282054423,0.003762675906796974,0.0037643381209897446,0.0037657791511514806,0.003766998806849806,0.003767996926888397,0.0037687733793375817,0.003769328061559401,0.003769660900227095,0.003769771851339039,0.003769660900227095,0.003769328061559401,0.0037687733793375817,0.003767996926888397,0.003766998806849806,0.0037657791511514806,0.0037643381209897446,0.003762675906796974,0.0037607927282054423,0.0037586888340056354,0.0037563645020990393,0.003753820039445428,0.003751055782004644,0.0037480720946729113,0.0037448693712136736,0.003741448034183014,0.0037378085348496225,0.003733951353109393,0.003729876997394628,0.0037255860045779,0.0037210789398705924,0.003716356396716135,0.0037114189966779842,0.003706267389322367,0.003700902252095814,0.003695324290197536,0.003689534236446657,0.0036835328511443557,0.0036773209219309456,0.003670899263637934,0.003664268718135102,0.0036574301541726453,0.0036503844672184198,0.003643132579290336,0.003635675438783951,0.003628014020295289,0.003620149324438965,0.0036120823776616346,0.0036038142320508415,0.0035953459651392886,0.0035866786797046145,0.0035778135035647017,0.0035687515893685936,0.0035594941143830563,0.0035500422802748535,0.0035403973128887893,0.0035305604620215728,0.0035205330011915718,0.003510316227404508,0.003499911460915155,0.003489320044985109,0.003478543345636684,0.003467582751403001,0.0034564396730743345,0.003445115543440783,0.0034336118170313202,0.0034219299698493052,0.0034100714991045097,0.0033980379229417317,0.003385830780166072,0.003373451629964919,0.0033609020516267457,0.003348183644256752,0.0033352980264894495,0.0033222468361982496,0.003309031730202117,0.0032956543839693835,0.0032821164913187538,0.003268419764117635,0.0032545659319777906,0.003240556741948457,0.0032263939582069497,0.0032120793617468574,0.0031976147500638874,0.0031830019368394302,0.0031682427516219382,0.003153339039506163,0.003138292660810352,0.003123105490751459,0.0031077794191184515,0.003092316349943788,0.0030767182011731393,0.003060986904333421,0.0030451244041992233,0.003029132658457702,0.0030130136373720065,0.0029967693234433175,0.0029804017110715746,0.0029639128062149554,0.0029473046260481885,0.0029305791986197725,0.002913738562508161,0.0028967847664770037,0.0028797198691295094,0.0028625459385619913,0.0028452650520166783,0.002827879295533866,0.0028103907636034633,0.002792801558816015,0.0027751137915132764,0.002757329579438388,0.0027394510473857424,0.002721480326850601,0.002703419555678523,0.002685270877714688,0.002667036442453171,0.0026487184046862303,0.0026303189241536954,0.002611840165192486,0.00259328429638637,0.0025746534902159855,0.0025559499227092173,0.002537175773091972,0.0025183332234394364,0.002499424458327856,0.0024804516644869132,0.0024614170304527666,0.0024423227462217895,0.002423171002905102,0.0024039639923839223,0.0023847039069658156,0.0023653929390418994,0.00234603328074504,0.0023266271236091285,0.002307176658229464,0.0022876840739243184,0.0022681515583977247,0.0022485812974035505,0.002228975474410903,0.0022093362702709273,0.0021896658628850364,0.00216996642687464,0.0021502401332524055,0.002130489149095115,0.0021107156372181584,0.0020909217558517205,0.0020711096583186915,0.0020512814927143696,0.002031439401587993,0.0020115855216261396,0.001991721983338051,0.001971850910742915,0.0019519744210591676,0.0019320946243958294,0.0019122136234459507,0.0018923335131821783,0.0018724563805545078,0.0018525843041902507,0.0018327193540962532,0.001812863591363419,0.00179301906787356,0.0017731878260086264,0.0017533718983623375,0.0017335733074542753,0.001713794065446446,0.0016940361738623725,0.0016743016233087364,0.0016545923931996142,0.0016349104514833332,0.0016152577543719858,0.0015956362460736399,0.0015760478585272663,0.001556494511140425,0.0015369781105297375,0.0015175005502641816,0.001498063710611228,0.0014786694582858606,0.0014593196462025088,0.00144001611322991,0.0014207606839489464,0.0014015551684134727,0.0013824013619141713,0.0013633010447454527,0.0013442559819754382,0.0013252679232190468,0.0013063386024142103,0.001287469737601248,0.0012686630307054232,0.0012499201673227068,0.001231242816508769,0.0012126326305712388,0.0011940912448652296,0.0011756202775921821,0.0011572213296020273,0.0011388959841987013,0.0011206458069490362,0.001102472345495047,0.0010843771293696303,0.0010663616698157123,0.0010484274596088495,0.0010305759728833177,0.0010128086649616977,9.951269721879936E-4,9.775323117642836E-4,9.600260815909479E-4,9.426096601104665E-4,9.25284406154831E-4,9.080516587965724E-4,8.909127372034287E-4,8.738689404966794E-4,8.569215476131493E-4,8.400718171709102E-4,8.233209873386998E-4,8.066702757090665E-4,7.901208791752656E-4,7.736739738119159E-4,7.573307147594434E-4,7.41092236112319E-4,7.249596508111086E-4,7.089340505383558E-4,6.930165056183088E-4,6.772080649205063E-4,6.61509755767235E-4,6.45922583844885E-4,6.304475331191992E-4,6.150855657544465E-4,5.998376220365209E-4,5.847046202999914E-4,5.69687456859102E-4,5.547870059427447E-4,5.400041196334158E-4,5.253396278101634E-4,5.10794338095539E-4,4.96369035806571E-4,4.820644839097579E-4,4.6788142298010544E-4,4.5382057116420525E-4,4.3988262414737674E-4,4.2606825512486865E-4,4.1237811477713975E-4,3.988128312492175E-4,3.8537301013415496E-4,3.720592344605779E-4,3.5887206468433925E-4,3.4581203868428665E-4,3.328796717621447E-4,3.2007545664651776E-4,3.0739986350102424E-4,2.9485333993655577E-4,2.82436311027678E-4,2.701491793331621E-4,2.5799232492066244E-4,2.4596610539553266E-4,2.340708559337868E-4,2.223068893192031E-4,2.1067449598457418E-4,1.9917394405709842E-4,1.8780547940791477E-4,1.7656932570577505E-4,1.6546568447485863E-4,1.544947351567141E-4,1.436566351763377E-4,1.3295152001236983E-4,1.2237950327141585E-4,1.1194067676647672E-4,1.0163511059948344E-4,9.146285324793341E-5,8.142393165561031E-5,7.151835132738339E-5,6.174609642807749E-5,5.210712988539563E-5,4.260139349688798E-5,3.322880804094929E-5,2.398927339183627E-5,1.4882668638683254E-5,5.9088522085035684E-6,-2.9323380068394464E-6,-1.1641084519710755E-5,-2.0217590111854238E-5,-2.866207769562532E-5,-3.697479017134127E-5,-4.51559902807569E-5,-5.320596045669486E-5,-6.112500266886022E-5,-6.891343826585312E-5,-7.657160781341133E-5,-8.409987092891577E-5,-9.149860611217436E-5,-9.876821057252495E-5,-1.0590910005228389E-4,-1.129217086465683E-4,-1.1980648861953246E-4,-1.2656391021704545E-4,-1.3319446147584584E-4,-1.3969864802921707E-4,-1.460769929092096E-4,-1.5233003634545404E-4,-1.5845833556061003E-4,-1.6446246456247804E-4,-1.7034301393283207E-4,-1.7610059061300354E-4,-1.8173581768626538E-4,-1.872493341570665E-4,-1.92641794727154E-4,-1.9791386956863696E-4,-2.030662440940416E-4,-2.0809961872340194E-4,-2.1301470864844454E-4,-2.178122435939148E-4,-2.2249296757609978E-4,-2.2705763865860155E-4,-2.3150702870542182E-4,-2.3584192313140493E-4,-2.4006312065010996E-4,-2.4417143301916003E-4,-2.481676847831353E-4,-2.520527130140718E-4,-2.558273670496255E-4,-2.594925082289659E-4,-2.6304900962646776E-4,-2.664977557832615E-4,-2.698396424367137E-4,-2.7307557624790357E-4,-2.76206474527165E-4,-2.792332649577624E-4,-2.82156885317778E-4,-2.849782832002719E-4,-2.8769841573179905E-4,-2.9031824928935014E-4,-2.9283875921579165E-4,-2.9526092953388724E-4,-2.9758575265896787E-4,-2.9981422911033533E-4,-3.0194736722147637E-4,-3.039861828491633E-4,-3.059316990815251E-4,-3.0778494594516987E-4,-3.095469601114339E-4,-3.1121878460185174E-4,-3.1280146849291723E-4,-3.142960666202276E-4,-3.1570363928209473E-4,-3.170252519427021E-4,-3.182619749349009E-4,-3.1941488316272813E-4,-3.2048505580373015E-4,-3.2147357601118576E-4,-3.2238153061631006E-4,-3.2321000983053124E-4,-3.2396010694792706E-4,-3.246329180479088E-4,-3.2522954169824546E-4,-3.2575107865851426E-4,-3.2619863158406774E-4,-3.2657330473060954E-4,-3.268762036594662E-4,-3.2710843494364805E-4,-3.2727110587478563E-4,-3.273653241710388E-4,-3.2739219768606074E-4,-3.273528341191147E-4,-3.272483407264294E-4,-3.270798240338866E-4,-3.268483895511276E-4,-3.265551414871733E-4,-3.2620118246764416E-4,-3.2578761325367155E-4,-3.2531553246258917E-4,-3.247860362904955E-4,-3.2420021823677324E-4,-3.235591688306561E-4,-3.2286397535993155E-4,-3.22115721601865E-4,-3.2131548755643383E-4,-3.2046434918195707E-4,-3.19563378133208E-4,-3.1861364150209177E-4,-3.1761620156097717E-4,-3.1657211550876086E-4,-3.1548243521975267E-4,-3.143482069954589E-4,-3.131704713193515E-4,-3.1195026261469406E-4,-3.1068860900551566E-4,-3.093865320808018E-4,-3.080450466619849E-4,-3.066651605738095E-4,-3.0524787441864803E-4,-3.037941813543404E-4,-3.0230506687563296E-4,-3.007815085992852E-4,-2.9922447605291937E-4,-2.976349304676783E-4,-2.960138245747612E-4,-2.943621024059075E-4,-2.9268069909788627E-4,-2.909705407010634E-4,-2.8923254399210543E-4,-2.8746761629087875E-4,-2.856766552816095E-4,-2.8386054883835577E-4,-2.82020174854853E-4,-2.8015640107878633E-4,-2.782700849505394E-4,-2.7636207344647806E-4,-2.7443320292681064E-4,-2.724842989880783E-4,-2.7051617632032027E-4,-2.6852963856895644E-4,-2.66525478201431E-4,-2.645044763786608E-4,-2.624674028313193E-4,-2.604150157410026E-4,-2.583480616263057E-4,-2.562672752338433E-4,-2.541733794342482E-4,-2.520670851231749E-4,-2.499490911273343E-4,-2.478200841155872E-4,-2.456807385151158E-4,-2.4353171643269812E-4,-2.4137366758110148E-4,-2.3920722921061115E-4,-2.370330260457115E-4,-2.3485167022692973E-4,-2.326637612578528E-4,-2.304698859573269E-4,-2.2827061841684395E-4,-2.2606651996312025E-4,-2.2385813912586836E-4,-2.2164601161076068E-4,-2.1943066027758476E-4,-2.172125951235829E-4,-2.1499231327196932E-4,-2.1277029896561763E-4,-2.1054702356590533E-4,-2.083229455567016E-4,-2.060985105534836E-4,-2.0387415131756386E-4,-2.0165028777540683E-4,-1.9942732704301277E-4,-1.9720566345534654E-4,-1.949856786007816E-4,-1.9276774136053326E-4,-1.9055220795304766E-4,-1.8833942198331612E-4,-1.861297144970781E-4,-1.839234040398753E-4,-1.8172079672091907E-4,-1.7952218628172918E-4,-1.773278541694991E-4,-1.751380696151447E-4,-1.729530897159882E-4,-1.707731595230259E-4,-1.6859851213273206E-4,-1.6642936878334233E-4,-1.6426593895556307E-4,-1.6210842047764885E-4,-1.5995699963478998E-4,-1.5781185128274774E-4,-1.556731389656764E-4,-1.5354101503806578E-4,-1.5141562079073928E-4,-1.492970865808406E-4,-1.4718553196573517E-4,-1.4508106584076137E-4,-1.4298378658075266E-4,-1.4089378218525974E-4,-1.3881113042739677E-4,-1.3673589900623043E-4,-1.346681457026374E-4,-1.326079185385475E-4,-1.3055525593948954E-4,-1.2851018690035904E-4,-1.2647273115432201E-4,-1.2444289934476804E-4,-1.224206932002273E-4,-1.204061057121627E-4,-1.1839912131554572E-4,-1.1639971607212963E-4,-1.1440785785632266E-4,-1.1242350654357457E-4,-1.1044661420117793E-4,-1.0847712528139286E-4,-1.065149768167974E-4,-1.0456009861776952E-4,-1.0261241347200124E-4,-1.0067183734594933E-4,-9.873827958812245E-5,-9.681164313410566E-5,-9.48918247132236E-5,-9.297871505674132E-5,-9.10721991075013E-5,-8.917215623089688E-5,-8.72784604270788E-5,-8.539098054429423E-5,-8.35095804932554E-5,-8.163411946243434E-5,-7.976445213418295E-5,-7.79004289015743E-5,-7.604189608586106E-5,-7.418869615445064E-5,-7.234066793929237E-5,-7.049764685557237E-5,-6.865946512061758E-5,-6.682595197290053E-5,-6.499693389104716E-5,-6.317223481274333E-5,-6.135167635343702E-5,-5.953507802473751E-5" />
-- Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
-- Retrieval info: 	<generic name="coeffScaling" value="Auto" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="8" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="Signed Binary" />
-- Retrieval info: 	<generic name="outMSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="18" />
-- Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
