-- megafunction wizard: %FIR Compiler II v13.1%
-- GENERATION: XML
-- LP100.vhd

-- Generated using ACDS version 13.1 162 at 2019.05.14.10:47:19

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LP100 is
	port (
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0';             --                     rst.reset_n
		ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(23 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0)                      --                        .error
	);
end entity LP100;

architecture rtl of LP100 is
	component LP100_0002 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(23 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component LP100_0002;

begin

	lp100_inst : component LP100_0002
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of LP100
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2019 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
-- Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
-- Retrieval info: 	<generic name="filterType" value="Single Rate" />
-- Retrieval info: 	<generic name="interpFactor" value="1" />
-- Retrieval info: 	<generic name="decimFactor" value="1" />
-- Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
-- Retrieval info: 	<generic name="clockRate" value="50" />
-- Retrieval info: 	<generic name="clockSlack" value="0" />
-- Retrieval info: 	<generic name="speedGrade" value="Medium" />
-- Retrieval info: 	<generic name="coeffReload" value="false" />
-- Retrieval info: 	<generic name="baseAddress" value="0" />
-- Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
-- Retrieval info: 	<generic name="backPressure" value="false" />
-- Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
-- Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
-- Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
-- Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
-- Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
-- Retrieval info: 	<generic name="inputRate" value="0.008" />
-- Retrieval info: 	<generic name="inputChannelNum" value="1" />
-- Retrieval info: 	<generic name="inputType" value="Signed Binary" />
-- Retrieval info: 	<generic name="inputBitWidth" value="24" />
-- Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="coeffSetRealValue" value="0.003585002057282315,0.0036209133948513724,0.0036841503417371553,0.0037744862631139604,0.003891487678530191,0.0040345215060500934,0.004202765277716284,0.004395220064380232,0.004610725783022638,0.0048479785046479625,0.00510554933732393,0.005381904428206455,0.005675425611281182,0.005984431224456947,0.006307196630495991,0.006641974000539617,0.0069870109557287775,0.007340567710269951,0.007700932416548395,0.008066434477542695,0.008435455661624012,0.008806438927464794,0.009177894939806914,0.009548406327842969,0.00991662980464612,0.010281296326326789,0.01064120952153652,0.010995242664036028,0.011342334492119415,0.011681484197967494,0.012011745917146965,0.01233222304356858,0.012642062678784345,0.01294045049746063,0.013226606274495683,0.013499780275155516,0.013759250659632719,0.014004321999622113,0.014234324948994185,0.014448617055596842,0.014646584648739157,0.014827645688985064,0.014991253425286025,0.015136900670713785,0.015264124483302437,0.015372511023590689,0.015461700355798602,0.01553139096519884,0.015581343779769273,0.01561138550887272,0.015621411144377194,0.01561138550887272,0.015581343779769273,0.01553139096519884,0.015461700355798602,0.015372511023590689,0.015264124483302437,0.015136900670713785,0.014991253425286025,0.014827645688985064,0.014646584648739157,0.014448617055596842,0.014234324948994185,0.014004321999622113,0.013759250659632719,0.013499780275155516,0.013226606274495683,0.01294045049746063,0.012642062678784345,0.01233222304356858,0.012011745917146965,0.011681484197967494,0.011342334492119415,0.010995242664036028,0.01064120952153652,0.010281296326326789,0.00991662980464612,0.009548406327842969,0.009177894939806914,0.008806438927464794,0.008435455661624012,0.008066434477542695,0.007700932416548395,0.007340567710269951,0.0069870109557287775,0.006641974000539617,0.006307196630495991,0.005984431224456947,0.005675425611281182,0.005381904428206455,0.00510554933732393,0.0048479785046479625,0.004610725783022638,0.004395220064380232,0.004202765277716284,0.0040345215060500934,0.003891487678530191,0.0037744862631139604,0.0036841503417371553,0.0036209133948513724,0.003585002057282315" />
-- Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
-- Retrieval info: 	<generic name="coeffScaling" value="Auto" />
-- Retrieval info: 	<generic name="coeffBitWidth" value="8" />
-- Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
-- Retrieval info: 	<generic name="outType" value="Signed Binary" />
-- Retrieval info: 	<generic name="outMSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outMsbBitRem" value="0" />
-- Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
-- Retrieval info: 	<generic name="outLsbBitRem" value="15" />
-- Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
-- Retrieval info: 	<generic name="bankCount" value="1" />
-- Retrieval info: 	<generic name="bankDisplay" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : NONE
